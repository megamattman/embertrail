library verilog;
use verilog.vl_types.all;
entity Embertrail_ctrl_vlg_tst is
end Embertrail_ctrl_vlg_tst;
